
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;
use ieee.math_real.all;
use std.textio.all;
use ieee.std_logic_textio.all;

package sim_file_pkg is
  ------------------------------------------------------------------------------
  -- Data Types
  ------------------------------------------------------------------------------
  type sim_file_bin_type            is file of character;

end sim_file_pkg;


package body sim_file_pkg is

end sim_file_pkg;