library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity maxMin is
generic(
  constant G_PIXEL_DEPTH   : integer := 16
);
Port();
end MaxMin;

architecture Behavioral of MaxMin is
begin